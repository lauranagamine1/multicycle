`timescale 1ns / 1ps

module HexTo7Segment (
    input wire [3:0] digit, 
    output reg [6:0] catode);
    
    always @(*) begin
        casex(digit) 
            4'b0000: catode = 7'b0111111; //0
            4'b0001: catode = 7'b0000110; //1
            4'b0010: catode = 7'b1011011; //2
            4'b0011: catode = 7'b1001111; //3
            4'b0100: catode = 7'b1100110; //4
            4'b0101: catode = 7'b1101101; //5
            4'b0110: catode = 7'b1111101; //6
            4'b0111: catode = 7'b0000111; //7
            4'b1000: catode = 7'b1111111; //8
            4'b1001: catode = 7'b1100111; //9
            4'b1010: catode = 7'b1110111; //A 
            4'b1011: catode = 7'b1111100; //B 
            4'b1100: catode = 7'b0111001; //C 
            4'b1101: catode = 7'b1011110; //D 
            4'b1110: catode = 7'b1111001; //E 
            4'b1111: catode = 7'b1110001; //F
            default: catode = 7'b0000000; // off
       endcase
    end
endmodule

module CLKdivider (
    input  wire        in_clk,
    input  wire        reset,    // reset asíncrono, activo alto
    output reg         out_clk
);

    // contador de 25 bits (genera un toggle cada vez que desborda)
    reg [24:0] counter;

    // reset asíncrono + lógica de división
    always @(posedge in_clk or posedge reset) begin
        if (reset) begin
            counter <= 0;
            out_clk <= 0;
        end else begin
            counter <= counter + 1;
            if (counter == 0)
                out_clk <= ~out_clk;
        end
    end

endmodule

module hFSM(input clk,input reset,input[15:0] data,output reg[3:0]
    digit,output reg[3:0] anode);
    
    reg [1:0] state;

    always @(posedge clk or posedge reset) begin
        if (reset)
            state <= 2'd0;
        else
            state <= state + 1'b1;
    end

    always @(*) begin
        case (state)
            2'd0: begin
                digit <= data[15:12];  // nibble más significativo
                anode <= 4'b0111;      // activa físicamente el dígito 3
            end
            2'd1: begin
                digit <= data[11: 8];
                anode <= 4'b1011;      // activa el dígito 2
            end
            2'd2: begin
                digit <= data[ 7: 4];
                anode <= 4'b1101;      // dígito 1
            end
            2'd3: begin
                digit <= data[ 3: 0];  // nibble menos significativo
                anode <= 4'b1110;      // dígito 0
            end
            default: begin
                digit <= 4'd0;
                anode <= 4'b1111;      // todos apagados
            end
        endcase
    end

endmodule

// Main module
module hex_display(input clk, input reset, input[15:0] data, output
    wire[3:0]anode, output wire[6:0]catode);
    wire scl_clk;
    wire[3:0] digit;
    CLKdivider sc(
        .in_clk(clk),
        .reset(reset),
        .out_clk(scl_clk)
    );
    hFSM m(
        .clk(scl_clk),
        .reset(reset),
        .data(data),
        .digit(digit),
        .anode(anode)
    );
    HexTo7Segment decoder (
        .digit(digit),
        .catode(catode)
    );
endmodule
